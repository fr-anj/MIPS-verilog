module ROM(
	input I_CLK,
	//input I_EN,
	
	input [7:0] I_ADDR,
	
	output reg [15:0] O_INSTR
);
	//internal variable or register declaration
	// N/A
	
	//implementation
	//clocked
	always @(posedge I_CLK) begin
		//if(I_EN) begin
			case(I_ADDR)
0: O_INSTR <= 16'b1100100100000000;
1: O_INSTR <= 16'b1100100000000010;
2: O_INSTR <= 16'b1101100101100111;
3: O_INSTR <= 16'b1010000101100111;
4: O_INSTR <= 16'b1011000111111000;


5: O_INSTR <= 16'b1100110100000000;
6: O_INSTR <= 16'b0010111010001001;
7: O_INSTR <= 16'b0011011110001001;
8: O_INSTR <= 16'b0011100010001111;
9: O_INSTR <= 16'b0100000110011001;
10: O_INSTR <= 16'b1100110000000000;
11: O_INSTR <= 16'b1100110111111111;
12: O_INSTR <= 16'b0101101011001101;
13: O_INSTR <= 16'b0110001011001101;
14: O_INSTR <= 16'b0110101011001101;
15: O_INSTR <= 16'b0111001011001101;
16: O_INSTR <= 16'b0111101011001101;
17: O_INSTR <= 16'b1000001011001101;
18: O_INSTR <= 16'b1100110011111111;
19: O_INSTR <= 16'b1100110100000000;
20: O_INSTR <= 16'b0101101011001101;
21: O_INSTR <= 16'b0110001011001101;
22: O_INSTR <= 16'b0110101011001101;
23: O_INSTR <= 16'b0111001011001101;
24: O_INSTR <= 16'b0111101011001101;
25: O_INSTR <= 16'b1000001011001101;
26: O_INSTR <= 16'b1100110000000000;
27: O_INSTR <= 16'b1100110111111111;
28: O_INSTR <= 16'b0101101011001101;
29: O_INSTR <= 16'b0110001011001101;
30: O_INSTR <= 16'b0110101011001101;
31: O_INSTR <= 16'b0111001011001101;
32: O_INSTR <= 16'b0111101011001101;
33: O_INSTR <= 16'b1000001011001101;
34: O_INSTR <= 16'b1100100010101010;
35: O_INSTR <= 16'b1100100100000011;
36: O_INSTR <= 16'b0001101010001001;
37: O_INSTR <= 16'b0010001010001001;
38: O_INSTR <= 16'b1100101110101010;
39: O_INSTR <= 16'b1100110010101010;
40: O_INSTR <= 16'b1100110100001000;
41: O_INSTR <= 16'b0001111011001101;
42: O_INSTR <= 16'b0010011011001101;
43: O_INSTR <= 16'b1100100000001111;
44: O_INSTR <= 16'b1100100100000100;
45: O_INSTR <= 16'b0001000010001001;
46: O_INSTR <= 16'b0000101010001001;
47: O_INSTR <= 16'b0000001010001001;
48: O_INSTR <= 16'b1100111000001111;
49: O_INSTR <= 16'b1100111111111111;
50: O_INSTR <= 16'b0100110111101111;
51: O_INSTR <= 16'b0101010111101111;
52: O_INSTR <= 16'b1000110111101111;
53: O_INSTR <= 16'b1100100000000000;
54: O_INSTR <= 16'b1100100100000000;
55: O_INSTR <= 16'b1100101000000000;
56: O_INSTR <= 16'b1100101100000000;
57: O_INSTR <= 16'b1101100000000000;
58: O_INSTR <= 16'b1101100100001111;
59: O_INSTR <= 16'b1101101011110000;
60: O_INSTR <= 16'b1101101111111111;
61: O_INSTR <= 16'b1100100001000011;
62: O_INSTR <= 16'b1101010000001111;
63: O_INSTR <= 16'b1101010100000000;
64: O_INSTR <= 16'b1101011011110000;
65: O_INSTR <= 16'b1101011111111111;
66: O_INSTR <= 16'b1100011111111000;
67: O_INSTR <= 16'b1100100001000110;
68: O_INSTR <= 16'b1101100000100011;
69: O_INSTR <= 16'b1011111100100011;
70: O_INSTR <= 16'b1100111111111111;
71: O_INSTR <= 16'b1100111001001101;
72: O_INSTR <= 16'b1101111001101001;
73: O_INSTR <= 16'b1100110111111111;
74: O_INSTR <= 16'b1001110101101001;
75: O_INSTR <= 16'b1100100000000000;
76: O_INSTR <= 16'b1100100100000000;
77: O_INSTR <= 16'b1100111000000000;
78: O_INSTR <= 16'b1101111001101001;
79: O_INSTR <= 16'b1100110100000000;
80: O_INSTR <= 16'b1001110101101001;
81: O_INSTR <= 16'b1100100001010110;
82: O_INSTR <= 16'b1101100001101001;
83: O_INSTR <= 16'b1100100100000000;
84: O_INSTR <= 16'b1010000101101001;
85: O_INSTR <= 16'b1100100011111111;
86: O_INSTR <= 16'b1100100000000000;
87: O_INSTR <= 16'b1101100001101001;
88: O_INSTR <= 16'b1100100100000001;
89: O_INSTR <= 16'b1010000101101001;
90: O_INSTR <= 16'b1100100000000000;
91: O_INSTR <= 16'b1101100001101001;
92: O_INSTR <= 16'b1100100100000000;
93: O_INSTR <= 16'b1010100111111000;
94: O_INSTR <= 16'b1100100001100011;
95: O_INSTR <= 16'b1101100001101001;
96: O_INSTR <= 16'b1100100111111111;
97: O_INSTR <= 16'b1010100111111000;
98: O_INSTR <= 16'b1100100000000000;
99: O_INSTR <= 16'b1100100000000000;
100: O_INSTR <= 16'b1101100001101001;
101: O_INSTR <= 16'b1100100111111111;
102: O_INSTR <= 16'b1011000111111000;
103: O_INSTR <= 16'b1100100001101101;
104: O_INSTR <= 16'b1101100001101001;
105: O_INSTR <= 16'b1100100100000000;
106: O_INSTR <= 16'b1011000111111000;
107: O_INSTR <= 16'b1100111100000000;
108: O_INSTR <= 16'b1100100000000000;
109: O_INSTR <= 16'b1100100100000000;
110: O_INSTR <= 16'b1100101000000000;
111: O_INSTR <= 16'b1100101100000000;
112: O_INSTR <= 16'b1100110000000000;
113: O_INSTR <= 16'b1100110100000000;
114: O_INSTR <= 16'b1100111000000000;
115: O_INSTR <= 16'b1100111100000000;
116: O_INSTR <= 16'b1100100000000000;
117: O_INSTR <= 16'b0010100110001000;
118: O_INSTR <= 16'b1100101000000000;
119: O_INSTR <= 16'b1100101100000000;
120: O_INSTR <= 16'b1100110000000000;
121: O_INSTR <= 16'b1100110100000000;
122: O_INSTR <= 16'b1100111000000000;
123: O_INSTR <= 16'b1100111100000000;
124: O_INSTR <= 16'b1100100000000000;
125: O_INSTR <= 16'b1100100100000000;
126: O_INSTR <= 16'b0010101010001000;
127: O_INSTR <= 16'b1100101100000000;
128: O_INSTR <= 16'b1100110000000000;
129: O_INSTR <= 16'b1100110100000000;
130: O_INSTR <= 16'b1100111000000000;
131: O_INSTR <= 16'b1100111100000000;
132: O_INSTR <= 16'b1100100000000000;
133: O_INSTR <= 16'b1100100100000000;
134: O_INSTR <= 16'b1100101000000000;
135: O_INSTR <= 16'b0010101110001000;
136: O_INSTR <= 16'b1100100000000000;
137: O_INSTR <= 16'b1100100100000000;
138: O_INSTR <= 16'b1100101000000000;
139: O_INSTR <= 16'b1100101100000000;
140: O_INSTR <= 16'b1100110000000000;
141: O_INSTR <= 16'b1100110100000000;
142: O_INSTR <= 16'b1100111000000000;
143: O_INSTR <= 16'b1100111100000000;
144: O_INSTR <= 16'b1100100010010110;
145: O_INSTR <= 16'b1111111111111111;
146: O_INSTR <= 16'b1111111111111111;
147: O_INSTR <= 16'b1111111111111111;
148: O_INSTR <= 16'b1111111111111111;
149: O_INSTR <= 16'b1111111111111111;
150: O_INSTR <= 16'b1100011111111000;


				default: O_INSTR <= 16'hFFFF;
			endcase
		//end
	end
	
endmodule 